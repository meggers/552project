module adder(in1, in2, out, control,  zr, neg);

input [15:0] in1, in2;
input [3:0] control;
output [15:0] out;
output zr, neg;
% output flags




endmodule
