module FU();

endmodule
