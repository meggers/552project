module cpu(clk, rst_n, hlt, pc);

//** DEFINE I/O INTERFACE **//
input clk;        	// Global clock signal
input rst_n;      	// Reset signal, active on low
output reg hlt;       	// Halt signal
output reg [15:0] pc; 	// Program counter

//** DEFINE GLOBAL VARS **//
localparam Z = 0;	// Index for Zero flag
localparam V = 1;	// Index for Overflow flag
localparam N = 2;	// Index for Sign flag

localparam RegWrite = 0;
localparam MemToReg = 1;
localparam MemWrite = 2;
localparam MemRead  = 3;
localparam PCSrc    = 4;
localparam ALUSrc   = 5;
localparam ALUOpLSB = 6;
localparam ALUOpMSB = 8;

localparam IF_ID_PC    = 0;
localparam IF_ID_INST  = 1;

localparam ID_EX_PC    = 0;
localparam ID_EX_OP1   = 1;
localparam ID_EX_OP2   = 2;
localparam ID_EX_INST  = 3;
localparam ID_EX_R0    = 0;
localparam ID_EX_R1    = 1;

localparam EX_MEM_PC   = 0;
localparam EX_MEM_RSLT = 1;
localparam EX_MEM_OP2  = 2;

localparam MEM_WB_RD   = 0;
localparam MEM_WB_RSLT = 1;

//** DEFINE REGISTERS **//
reg [2:0] FLAG;		// Flag register

reg [8:0] CTRL_ID_EX;
reg [4:0] CTRL_EX_MEM;
reg [1:0] CTRL_MEM_WB;

reg [15:0] DATA_IF_ID [1:0];
reg [15:0] DATA_ID_EX [3:0];
reg [15:0] DATA_EX_MEM [2:0];
reg [15:0] DATA_MEM_WB [1:0];

reg [3:0] REG_ID_EX [1:0];
reg [3:0] REG_EX_MEM;
reg [3:0] REG_MEM_WB;

//** DEFINE WIRES **//
wire [15:0] pc_incr, instr, read_1, 
	    read_2, dm_read, op_2,
	    result;

wire [8:0] ctrl_signals;

wire [2:0] flags;

//** DEFINE MODULES **//
IM instr_mem(.clk(clk), 		// INSTRUCTION MEMORY
	     .addr(pc), 
             .rd_en(),// TODO
	     .instr(instr));	
			
DM  data_mem(.clk(clk),			// DATA MEMORY
	     .addr(DATA_EX_MEM[EX_MEM_RSLT]),
	     .re(CTRL_EX_MEM[MemRead]), 
             .we(CTRL_EX_MEM[MemWrite]),
	     .wrt_data(DATA_EX_MEM[EX_MEM_OP2]),
	     .rd_data(dm_read));// TODO

rf  reg_file(.clk(clk), 		// REGISTER FILE
	     .p0_addr(DATA_IF_ID[IF_ID_INST][11:8]), 
	     .p1_addr(DATA_IF_ID[IF_ID_INST][7:4]), 
	     .p0(read_1), 
	     .p1(read_2),
	     .re0(), .re1(),// TODO 
	     .dst_addr(REG_MEM_WB), 
	     .dst(),// TODO 
	     .we(CTRL_MEM_WB[RegWrite]), 
	     .hlt(hlt));

Control ctrl(.instr(DATA_IF_ID[IF_ID_INST][15:12]),	// CONTROL BLOCK
	     .ctrl_signals(ctrl_signals));


module alu(.ALUop(CTRL_ID_EX[ALUOpMSB, ALUOpLSB]), 
	   .src0(DATA_ID_EX[ID_EX_OP1]), 
	   .src1(op_2), 
	   .result(result), 
	   .flags(flags));

//** CONTINUOUS ASSIGNS **//
assign pc_incr = pc + 4;
assign op_2 = CTRL_ID_EX[ALUSrc] ? {12'h000, DATA_ID_EX[ID_EX_INST][3:0]} : DATA_ID_EX[ID_EX_OP1];

//** PROGRAM COUNTER **//
always @(posedge clk or negedge rst_n) begin 
	if (~rst_n) begin
		pc <= 0;
	end else begin
		pc <= (CTRL_EX_MEM[PCSrc] & FLAG[Z]) ? DATA_EX_EM[EX_MEM_PC] : pc_incr;
	end
end

//** CONTROL PIPELINE **//
always @(posedge clk or negedge rst_n) begin
	if (~rst_n) begin
		CTRL_ID_EX  <= 0;
		CTRL_EM_MEM <= 0;
		CTRL_MEM_WB <= 0;
	end else begin
		CTRL_ID_EX  <= ctrl_signals;
		CTRL_EM_MEM <= CTRL_ID_EX[Branch:MemWrite];
		CTRL_MEM_WB <= CTRL_EM_MEM[MemToReg:RegWrite];
	end
end

//** DATA PIPELINE **//
always @(posedge clk or negedge rst_n) begin
	if (~rst_n) begin
		DATA_IF_ID <= 0; // TODO: this doesn't work
		DATA_ID_EX <= 0;
		DATA_EX_MEM <= 0;
		DATA_MEM_WB <= 0;
	end else begin
		DATA_IF_ID[IF_ID_PC] <= pc_incr;
		DATA_IF_ID[IF_ID_INST] <= instr;

		DATA_ID_EX[ID_EX_PC] <= DATA_IF_ID[IF_ID_PC];
		DATA_ID_EX[ID_EX_OP1] <= read_1;
		DATA_ID_EX[ID_EX_OP2] <= read_2;
		DATA_ID_EX[ID_EX_INST] <= DATA_IF_ID[IF_ID_INST];

		DATA_EX_MEM[EX_MEM_PC] <= DATA_ID_EX[ID_EX_PC];
		DATA_EX_MEM[EX_MEM_RSLT] <= result;
		FLAG <= flags;
		DATA_EX_MEM[EX_MEM_OP2] <= DATA_ID_EX[ID_EX_OP2];
		REG_EX_MEM <= DATA_ID_EX[ID_EX_INST][11:8];

		DATA_MEM_WB[MEM_WB_RD] <= dm_read;
		DATA_MEM_WB[MEM_WB_RSLT] <= DATA_EX_MEM[EX_MEM_RSLT];
		REG_MEM_WB <= REG_EX_MEM;
	end
end

module


endmodule Control(instr, ctrl_signals);

input [3:0] instr;
output [8:0] ctrl_signals;

localparam RegWrite = 0;
localparam MemToReg = 1;
localparam MemWrite = 2;
localparam MemRead  = 3;
localparam PCSrc    = 4;
localparam ALUSrc   = 5;
localparam RegDst   = 6;
localparam ALUOpLSB = 7;
localparam ALUUpMSB = 8;

endmodule


module aluControl(ALUOp, instr);

endmodule
