module HDU(instr, write_data, mem_read, pc_write, if_id_write, stall);

input [15:0] instr, write_data;
input mem_read;
output pc_write, if_id_write, stall;

endmodule
